* First line
.include "2um_CMOS.modlib"


*Definici�n de subcircuitos

* Inversor de 1w de dimension sin capacitancias parasitas
.subckt inv_1w_nopara nin nout nsup ngnd
Mpmos nout nin nsup nsup P_2u L=2u W=6u AD=36p PD=24u AS=36p PS=24u ;
Mnmos nout nin ngnd ngnd N_2u L=2u W=6u AD=36p PD=24u AS=36p PS=24u ;
.ends

* Inversor de 3w de dimension sin capacitancias parasitas
.subckt inv_3w_nopara nin nout nsup ngnd
Mpmos nout nin nsup nsup P_2u L=2u W=18u AD=108p PD=48u AS=108p PS=48u ;
Mnmos nout nin ngnd ngnd N_2u L=2u W=18u AD=108p PD=48u AS=108p PS=48u ;
.ends

* Inversor de 1w de dimension con capacitancias parasitas
.subckt inv_1w_para nin nout nsup ngnd
Mpmos nout nin nsup nsup P_2u L=2u W=6u AD=36p PD=24u AS=36p PS=24u ;
Mnmos nout nin ngnd ngnd N_2u L=2u W=6u AD=36p PD=24u AS=36p PS=24u ;

Cpar1 nsup 0 171.56183f
Cpar2 ngnd 0 137.77681f
Cpar3 nout 0 138.46099f
Cpar4 nin 0 8.9924632f
.ends

* Inversor de 3w de dimension con capacitancias parasitas
.subckt inv_3w_para nin nout nsup ngnd
Mpmos nout nin nsup nsup P_2u L=2u W=18u AD=108p PD=48u AS=108p PS=48u ;
Mnmos nout nin ngnd ngnd N_2u L=2u W=18u AD=108p PD=48u AS=108p PS=48u ;

Cpar1 nsup 0 472.94321f
Cpar2 ngnd 0 413.9192f
Cpar3 nout 0 412.03771f
Cpar4 nin 0 13.195057f
.ends


*Instanciamiento de circuiteria

* Inversor de 1w de dimension sin capacitancias parasitas
X_inv1w_nopara Vin vout_1w_nopara Vdd 0 inv_1w_nopara
X_inv3w_nopara Vin vout_3w_nopara Vdd 0 inv_3w_nopara
X_inv1w_para Vin vout_1w_para Vdd 0 inv_1w_para
X_inv3w_para Vin vout_3w_para Vdd 0 inv_3w_para

* Definici�n de Voltajes
Vdd Vdd 0 DC 5
Vin Vin 0 PULSE(5 0 0.01m 1p 1p 0.01m 0.02m 1)


*Definici�n de analisis
.tran 30u uic


* Analisis de dimensiones
* tp_LH
* 1w = 10.000262 us - 10 us
* 3w = 10.000248 us - 10 us

* tp_HL
* 1w = 20.000078 us - 20 us
* 3w = 20.000074 us - 20 us

* tp
* 1w = (262 ps + 78 ps )/2 = 170 ps
* 3w = (248 ps + 74 ps )/2 = 161 ps

* diferencia de tp
* 1w - 3w = 170 ps - 161 ps = 9 ps

* Analisis de parasitos

* 1w
* tp_LH
* para =    10.001156 us - 10 us
* no_para = 10.000262 us - 10 us

*tp_HL
* para =    20.000358 us - 20 us
* no_para = 20.000078 us - 20 us

*tp
* para =    (1156 ps + 358 ps )/2 = 757 ps
* no_para = (262 ps  + 78 ps  )/2 = 170 ps

*3w
* tp_LH
* para =    10.001122 us - 10 us
* no_para = 10.000248 us - 10 us

*tp_HL
* para =    20.000349 us - 20 us
* no_para = 20.000074 us - 20 us

*tp
* para =    (1122 ps + 349 ps )/2 = 735.5 ps
* no_para = (248 ps  + 74 ps  )/2 = 161 ps

